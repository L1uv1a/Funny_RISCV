module forward_tb (
);
    
endmodule